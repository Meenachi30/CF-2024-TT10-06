
`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.02.2025 21:23:07
// Design Name: 
// Module Name: clock_div
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module clock_div(
    input clk,        // Input clock (assumed 100 MHz for this example)
    input reset,         // Synchronous reset
    output reg w_clk,   // 50 MHz write clock output
    output reg r_clk    // 30 MHz read clock output
);

    reg [2:0] wr_counter = 3'b000;  // Counter for write clock division
    reg [2:0] rd_counter = 3'b000; // Counter for read clock division

    // Generate 50 MHz clock (divide by 1.2)
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            wr_counter <= 3'b000;
            w_clk <= 1'b0;
        end else if (wr_counter == 1) begin
            wr_counter <= 3'b000;
            w_clk <= ~w_clk;
        end else begin
            wr_counter <= wr_counter + 1'b1;
        end
    end

    // Generate 30 MHz clock (approximate divide by 2)
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            rd_counter <= 3'b000;
            r_clk <= 1'b0;
        end else if (rd_counter == 2) begin
            rd_counter <= 3'b000;
            r_clk <= ~r_clk;
        end else begin
            rd_counter <= rd_counter + 1'b1;
        end
    end



endmodule
